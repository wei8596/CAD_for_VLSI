module io(O,in,clk);

input clk;
input [7:0] in;

output [7:0] O;


assign O=in;




endmodule