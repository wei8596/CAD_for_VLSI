module test(O,clk);

input clk;


output [7:0] O;


assign O=~(8'b11110000);




endmodule